module comparator
#
(N = 8)
(
    input i_val,
    input [N-1:0] ref_high,
    input [N-1:0] ref_low,
    output o_fault
);

    assign o_fault = ;

endmodule
